** Profile: "SCHEMATIC1-transient"  [ C:\Users\razvan.cacu\Desktop\CAD\proiect\PROIECT CAD-PSpiceFiles\SCHEMATIC1\transient.sim ] 

** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\razvan.cacu\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\Users\razvan.cacu\Desktop\OPA847_MODEL.OLB" 
.lib "C:\Users\razvan.cacu\Desktop\CAD\lab7\ex1-PSpiceFiles\SCHEMATIC1\SCHEMATIC1.LIB" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 6ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
