** Profile: "SCHEMATIC1-monte carlo"  [ c:\users\razvan.cacu\desktop\proiect cad\cad-pspicefiles\schematic1\monte carlo.sim ] 

** Creating circuit file "monte carlo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 
.MC 20 TRAN v([OUT_TRI]) YMAX OUTPUT ALL SEED=400 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
